library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY mapping_tb is
END mapping_tb;

ARCHITECTURE Behavioral of mapping_tb is
begin

end ARCHITECTURE
